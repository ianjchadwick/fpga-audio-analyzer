`timescale 1ns / 1ps

// Generate HS, VS signals from pixel clock.
// hcounter & vcounter are the index of the current pixel 
// origin (0, 0) at top-left corner of the screen
// valid display range for hcounter: [0, 640)
// valid display range for vcounter: [0, 480)
module vga_controller_640_60 (pixel_clk,HS,VS,hcounter,vcounter,blank);

	input pixel_clk;
	output HS, VS, blank;
	output [10:0] hcounter, vcounter;

	parameter HMAX = 800; // maximum value for the horizontal pixel counter
	parameter VMAX = 525; // maximum value for the vertical pixel counter
	parameter HLINES = 640; // total number of visible columns
	parameter HFP = 648; // value for the horizontal counter where front porch ends
	parameter HSP = 744; // value for the horizontal counter where the synch pulse ends
	parameter VLINES = 480; // total number of visible lines
	parameter VFP = 482; // value for the vertical counter where the front porch ends
	parameter VSP = 484; // value for the vertical counter where the synch pulse ends
	parameter SPP = 0;


	wire video_enable;
	reg HS,VS,blank;
	reg [10:0] hcounter,vcounter;

	always@(posedge pixel_clk)begin
		blank <= ~video_enable; 
	end

	always@(posedge pixel_clk)begin
		if (hcounter == HMAX) hcounter <= 0;
		else hcounter <= hcounter + 1;
	end

	always@(posedge pixel_clk)begin
		if(hcounter == HMAX) begin
			if(vcounter == VMAX) vcounter <= 0;
			else vcounter <= vcounter + 1; 
		end
	end

	always@(posedge pixel_clk)begin
		if(hcounter >= HFP && hcounter < HSP) HS <= SPP;
		else HS <= ~SPP; 
	end

	always@(posedge pixel_clk)begin
		if(vcounter >= VFP && vcounter < VSP) VS <= SPP;
		else VS <= ~SPP; 
	end

	assign video_enable = (hcounter < HLINES && vcounter < VLINES) ? 1'b1 : 1'b0;

endmodule


// top module that instantiate the VGA controller and generate images
module vga_top(
    input clk,
    input [3:0] score,
    output reg [3:0] VGA_R,
    output reg [3:0] VGA_G,
    output reg [3:0] VGA_B,
    output wire VGA_HS,
    output wire VGA_VS
    );
    
localparam

R_BG = 4'h2,
G_BG = 4'h2,
B_BG = 4'h2,

SCORE_R_OFF = 4'h8,
SCORE_G_OFF = 4'h8,
SCORE_B_OFF = 4'h8,

SCORE_R_ON = 4'h0,
SCORE_G_ON = 4'h0,
SCORE_B_ON = 4'h0,

TOP_R_ON = 4'hF,
TOP_G_ON = 4'hF,
TOP_B_ON = 4'h3,

TOP_R_OFF = R_BG,
TOP_G_OFF = G_BG,
TOP_B_OFF = B_BG,

BOT_R_ON = 4'h6,
BOT_G_ON = 4'h0,
BOT_B_ON = 4'h6,

BOT_R_OFF = R_BG,
BOT_G_OFF = G_BG,
BOT_B_OFF = B_BG;


reg pclk_div_cnt;
reg pixel_clk;
reg [3:0] row_counter = 4'd0;
wire [10:0] vga_hcnt, vga_vcnt;
wire vga_blank;

reg [15:0] row0 = 16'd0,
           row1 = 16'd0,
           row2 = 16'd0,
           row3 = 16'd0,
           row4 = 16'd0,
           row5 = 16'd0,
           row6 = 16'd0,
           row7 = 16'd0,
           row8 = 16'd0,
           row9 = 16'd0,
           row10 = 16'd0,
           row11 = 16'd0,
           row12 = 16'd0,
           row13 = 16'd0,
           row14 = 16'd0,
           row15 = 16'd0;
           
           //"SCORE:"      
reg [47:0] top_row0  = 48'd0,
           top_row1  = 48'd0,
           top_row2  = {8'b01111100,8'b00111100,8'b01111100,8'b11111100,8'b11111110,8'b00000000},
           top_row3  = {8'b11000110,8'b01100110,8'b11000110,8'b01100110,8'b01100110,8'b00000000},
           top_row4  = {8'b11000110,8'b11000010,8'b11000110,8'b01100110,8'b01100010,8'b00011000},
           top_row5  = {8'b01100000,8'b11000000,8'b11000110,8'b01100110,8'b01101000,8'b00011000},
           top_row6  = {8'b00111000,8'b11000000,8'b11000110,8'b01111100,8'b01111000,8'b00000000},
           top_row7  = {8'b00001100,8'b11000000,8'b11000110,8'b01101100,8'b01101000,8'b00000000},
           top_row8  = {8'b00000110,8'b11000000,8'b11000110,8'b01100110,8'b01100000,8'b00000000},
           top_row9  = {8'b11000110,8'b11000010,8'b11000110,8'b01100110,8'b01100010,8'b00011000},
           top_row10 = {8'b11000110,8'b01100110,8'b11000110,8'b01100110,8'b01100110,8'b00011000},
           top_row11 = {8'b01111100,8'b00111100,8'b01111100,8'b11100110,8'b11111110,8'b00000000},
           top_row12 = 48'd0,
           top_row13 = 48'd0,
           top_row14 = 48'd0,
           top_row15 = 48'd0;                 
 
            //{music note}Krazy Karaoke!{music note}                
 reg [127:0] bot_row0  = {128'd0},
            bot_row1  = {128'd0},
            bot_row2  = {8'b00111111,8'b01100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11100000,8'b00000000,8'b00011000,8'b01111111},
            bot_row3  = {8'b00110011,8'b01100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b01100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b01100000,8'b00000000,8'b00111100,8'b01100011},
            bot_row4  = {8'b00111111,8'b01100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b01100110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b01100000,8'b00000000,8'b00111100,8'b01111111},
            bot_row5  = {8'b00110000,8'b01101100,8'b11011100,8'b01111000,8'b11111110,8'b11000110,8'b00000000,8'b01101100,8'b01111000,8'b11011100,8'b01111000,8'b01111100,8'b01100110,8'b01111100,8'b00111100,8'b01100011},
            bot_row6  = {8'b00110000,8'b01111000,8'b01110110,8'b00001100,8'b11001100,8'b11000110,8'b00000000,8'b01111000,8'b00001100,8'b01110110,8'b00001100,8'b11000110,8'b01101100,8'b11000110,8'b00011000,8'b01100011},
            bot_row7  = {8'b00110000,8'b01111000,8'b01100110,8'b01111100,8'b00011000,8'b11000110,8'b00000000,8'b01111000,8'b01111100,8'b01100110,8'b01111100,8'b11000110,8'b01111000,8'b11111110,8'b00011000,8'b01100011},
            bot_row8  = {8'b00110000,8'b01101100,8'b01100000,8'b11001100,8'b00110000,8'b11000110,8'b00000000,8'b01101100,8'b11001100,8'b01100000,8'b11001100,8'b11000110,8'b01111000,8'b11000000,8'b00011000,8'b01100011},
            bot_row9  = {8'b00110000,8'b01100110,8'b01100000,8'b11001100,8'b00110000,8'b11000110,8'b00000000,8'b01100110,8'b11001100,8'b01100000,8'b11001100,8'b11000110,8'b01101100,8'b11000000,8'b00000000,8'b01100111},
            bot_row10 = {8'b11110000,8'b01100110,8'b01100000,8'b11001100,8'b11000110,8'b11000110,8'b00000000,8'b01100110,8'b11001100,8'b01100000,8'b11001100,8'b11000110,8'b01100110,8'b11000110,8'b00011000,8'b11100111},
            bot_row11 = {8'b11100000,8'b11100110,8'b11110000,8'b01110110,8'b11111110,8'b01111110,8'b00000000,8'b11100110,8'b01110110,8'b11110000,8'b01110110,8'b01111100,8'b11100110,8'b01111100,8'b00011000,8'b11100110},
            bot_row12 = {8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000110,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11000000},
            bot_row13 = {8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00001100,8'b00000000,72'd0},
            bot_row14 = {8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b11111000,8'b00000000,72'd0},
            bot_row15 = {8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,72'd0};                

//Bits with a 1 are black 0 are white in the 320x320 grid in the center
//each case corresponds to displaying that digit
always@(score)begin
    case(score)
    4'd10:  begin
                 row0  = 16'b0000000000000000;
                 row1  = 16'b0000000000000000;
                 row2  = 16'b0001100001111100;
                 row3  = 16'b0011100011000110;
                 row4  = 16'b0111100011000110;
                 row5  = 16'b0001100011001110;
                 row6  = 16'b0001100011011110;
                 row7  = 16'b0001100011110110;
                 row8  = 16'b0001100011100110;
                 row9  = 16'b0001100011000110;
                 row10 = 16'b0001100011000110;
                 row11 = 16'b0111111001111100;
                 row12 = 16'b0000000000000000;
                 row13 = 16'b0000000000000000;
                 row14 = 16'b0000000000000000;
                 row15 = 16'b0000000000000000;
            end
    
    4'd9:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_01111100_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_11000110_0000;
                 row5  = 16'b0000_11000110_0000;
                 row6  = 16'b0000_01111110_0000;
                 row7  = 16'b0000_00000110_0000;
                 row8  = 16'b0000_00000110_0000;
                 row9  = 16'b0000_00000110_0000;
                 row10 = 16'b0000_00001100_0000;
                 row11 = 16'b0000_01111000_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    4'd8:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_01111100_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_11000110_0000;
                 row5  = 16'b0000_11000110_0000;
                 row6  = 16'b0000_01111100_0000;
                 row7  = 16'b0000_11000110_0000;
                 row8  = 16'b0000_11000110_0000;
                 row9  = 16'b0000_11000110_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_01111100_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    
    4'd7:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_11111110_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_00000110_0000;
                 row5  = 16'b0000_00000110_0000;
                 row6  = 16'b0000_00001100_0000;
                 row7  = 16'b0000_00011000_0000;
                 row8  = 16'b0000_00110000_0000;
                 row9  = 16'b0000_00110000_0000;
                 row10 = 16'b0000_00110000_0000;
                 row11 = 16'b0000_00110000_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
            
    4'd6:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_00111000_0000;
                 row3  = 16'b0000_01100000_0000;
                 row4  = 16'b0000_11000000_0000;
                 row5  = 16'b0000_11000000_0000;
                 row6  = 16'b0000_11111100_0000;
                 row7  = 16'b0000_11000110_0000;
                 row8  = 16'b0000_11000110_0000;
                 row9  = 16'b0000_11000110_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_01111100_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
            
    4'd5:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_11111110_0000;
                 row3  = 16'b0000_11000000_0000;
                 row4  = 16'b0000_11000000_0000;
                 row5  = 16'b0000_11000000_0000;
                 row6  = 16'b0000_11111100_0000;
                 row7  = 16'b0000_00000110_0000;
                 row8  = 16'b0000_00000110_0000;
                 row9  = 16'b0000_00000110_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_01111100_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
            
    4'd4:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_00001100_0000;
                 row3  = 16'b0000_00011100_0000;
                 row4  = 16'b0000_00111100_0000;
                 row5  = 16'b0000_01101100_0000;
                 row6  = 16'b0000_11001100_0000;
                 row7  = 16'b0000_11111110_0000;
                 row8  = 16'b0000_00001100_0000;
                 row9  = 16'b0000_00001100_0000;
                 row10 = 16'b0000_00001100_0000;
                 row11 = 16'b0000_00011110_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    
    4'd3:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_01111100_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_00000110_0000;
                 row5  = 16'b0000_00000110_0000;
                 row6  = 16'b0000_00111100_0000;
                 row7  = 16'b0000_00000110_0000;
                 row8  = 16'b0000_00000110_0000;
                 row9  = 16'b0000_00000110_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_01111100_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    
    4'd2:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_01111100_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_00000110_0000;
                 row5  = 16'b0000_00001100_0000;
                 row6  = 16'b0000_00011000_0000;
                 row7  = 16'b0000_00110000_0000;
                 row8  = 16'b0000_01100000_0000;
                 row9  = 16'b0000_11000000_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_11111110_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    
    4'd1:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_00011000_0000;
                 row3  = 16'b0000_00111000_0000;
                 row4  = 16'b0000_01111000_0000;
                 row5  = 16'b0000_00011000_0000;
                 row6  = 16'b0000_00011000_0000;
                 row7  = 16'b0000_00011000_0000;
                 row8  = 16'b0000_00011000_0000;
                 row9  = 16'b0000_00011000_0000;
                 row10 = 16'b0000_00011000_0000;
                 row11 = 16'b0000_01111110_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
            
    4'd0:   begin
                 row0  = 16'b0000_00000000_0000;
                 row1  = 16'b0000_00000000_0000;
                 row2  = 16'b0000_01111100_0000;
                 row3  = 16'b0000_11000110_0000;
                 row4  = 16'b0000_11000110_0000;
                 row5  = 16'b0000_11001110_0000;
                 row6  = 16'b0000_11011110_0000;
                 row7  = 16'b0000_11110110_0000;
                 row8  = 16'b0000_11100110_0000;
                 row9  = 16'b0000_11000110_0000;
                 row10 = 16'b0000_11000110_0000;
                 row11 = 16'b0000_01111100_0000;
                 row12 = 16'b0000_00000000_0000;
                 row13 = 16'b0000_00000000_0000;
                 row14 = 16'b0000_00000000_0000;
                 row15 = 16'b0000_00000000_0000;
            end
    
    default begin
                 row0 = 16'd0;
                 row1 = 16'd0;
                 row2 = 16'd0;
                 row3 = 16'd0;
                 row4 = 16'd0;
                 row5 = 16'd0;
                 row6 = 16'd0;
                 row7 = 16'd0;
                 row8 = 16'd0;
                 row9 = 16'd0;
                 row10 = 16'd0;
                 row11 = 16'd0;
                 row12 = 16'd0;
                 row13 = 16'd0;
                 row14 = 16'd0;
                 row15 = 16'd0;
            end
    
    endcase

end









// Clock divider. Generate 25MHz pixel_clk from 100MHz clock.
always @(posedge clk) begin
    pclk_div_cnt <= !pclk_div_cnt;
    if (pclk_div_cnt == 1'b1) pixel_clk <= !pixel_clk;
end



// Instantiate VGA controller
vga_controller_640_60 vga_controller(
    .pixel_clk(pixel_clk),
    .HS(VGA_HS),
    .VS(VGA_VS),
    .hcounter(vga_hcnt),
    .vcounter(vga_vcnt),
    .blank(vga_blank)
);

// Generate figure to be displayed
// Decide the color for the current pixel at index (hcnt, vcnt).
// This example displays an white square at the center of the screen with a colored checkerboard background.
always @(*) begin
    // Set pixels to black during Sync. Failure to do so will result in dimmed colors or black screens.
    if (vga_blank) begin 
        VGA_R = 0;
        VGA_G = 0;
        VGA_B = 0;
    end
    else begin  // Image to be displayed
        VGA_R = 4'h2;
        VGA_G = 4'h2;
        VGA_B = 4'h2;
        
        
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 1) && (vga_vcnt <= 5) ) ) begin
            if(top_row0[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 6) && (vga_vcnt <= 10) ) ) begin
            if(top_row1[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 11) && (vga_vcnt <= 15) ) ) begin
            if(top_row2[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 16) && (vga_vcnt <= 20) ) ) begin
            if(top_row3[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 21) && (vga_vcnt <= 25) ) ) begin
            if(top_row4[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 26) && (vga_vcnt <= 30) ) ) begin
            if(top_row5[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 31) && (vga_vcnt <= 35) ) ) begin
            if(top_row6[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 36) && (vga_vcnt <= 40) ) ) begin
            if(top_row7[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 41) && (vga_vcnt <= 45) ) ) begin
            if(top_row8[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 46) && (vga_vcnt <= 50) ) ) begin
            if(top_row9[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 51) && (vga_vcnt <= 55) ) ) begin
            if(top_row10[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 56) && (vga_vcnt <= 60) ) ) begin
            if(top_row11[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 61) && (vga_vcnt <= 65) ) ) begin
            if(top_row12[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 66) && (vga_vcnt <= 70) ) ) begin
            if(top_row13[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 71) && (vga_vcnt <= 75) ) ) begin
            if(top_row14[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[47] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[46] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[45] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[44] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[43] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[42] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[41] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[40] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[39] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[38] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[37] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[36] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[35] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[34] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[33] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[32] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[31] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[30] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[29] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[28] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[27] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[26] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[25] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[24] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[23] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[22] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[21] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[20] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[19] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[18] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[17] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[16] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[15] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[14] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[13] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[12] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[11] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[10] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[9] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[8] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[7] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[6] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[5] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[4] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[3] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[2] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[1] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 76) && (vga_vcnt <= 80) ) ) begin
            if(top_row15[0] == 1'b1)
                begin
                    VGA_R = TOP_R_ON;
                    VGA_G = TOP_G_ON;
                    VGA_B = TOP_B_ON;
                end
            else
                begin
                    VGA_R = TOP_R_OFF;
                    VGA_G = TOP_G_OFF;
                    VGA_B = TOP_B_OFF;
                end
            
            end
            

        /*************************SCORE SECTION******************************/
        
        //Centered 320x320 square matrix in 20x20 blocks [Row, Col]
        //Row0
        //[0,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
            if(row0[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[0,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 81 && vga_vcnt <= 100)) begin
			if(row0[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW1
        //[1,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[1,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 101 && vga_vcnt <= 120)) begin
			if(row1[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW2
        //[2,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[2,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 121 && vga_vcnt <= 140)) begin
			if(row2[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW3
        //[3,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[3,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 141 && vga_vcnt <= 160)) begin
			if(row3[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW4
        //[4,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[4,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 161 && vga_vcnt <= 180)) begin
			if(row4[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW5
        //[5,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[5,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 181 && vga_vcnt <= 200)) begin
			if(row5[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW6
        //[6,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[6,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 201 && vga_vcnt <= 220)) begin
			if(row6[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW7
        //[7,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[7,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 221 && vga_vcnt <= 240)) begin
			if(row7[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW8
        //[8,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[8,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 241 && vga_vcnt <= 260)) begin
			if(row8[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW9
        //[9,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[9,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 261 && vga_vcnt <= 280)) begin
			if(row9[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW10
        //[10,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[10,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 281 && vga_vcnt <= 300)) begin
			if(row10[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW11
        //[11,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[11,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 301 && vga_vcnt <= 320)) begin
			if(row11[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW12
        //[12,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[12,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 321 && vga_vcnt <= 340)) begin
			if(row12[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW13
        //[13,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[13,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 341 && vga_vcnt <= 360)) begin
			if(row13[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW14
        //[14,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[14,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 361 && vga_vcnt <= 380)) begin
			if(row14[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //ROW15
        //[15,0]
        if ((vga_hcnt >= 161 && vga_hcnt <= 180) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[15] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,1]
        if ((vga_hcnt >= 181 && vga_hcnt <= 200) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[14] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,2]
        if ((vga_hcnt >= 201 && vga_hcnt <= 220) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[13] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,3]
        if ((vga_hcnt >= 221 && vga_hcnt <= 240) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[12] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,4]
        if ((vga_hcnt >= 241 && vga_hcnt <= 260) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[11] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,5]
        if ((vga_hcnt >= 261 && vga_hcnt <= 280) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[10] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,6]
        if ((vga_hcnt >= 281 && vga_hcnt <= 300) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[9] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,7]
        if ((vga_hcnt >= 301 && vga_hcnt <= 320) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[8] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,8]
        if ((vga_hcnt >= 321 && vga_hcnt <= 340) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[7] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,9]
        if ((vga_hcnt >= 341 && vga_hcnt <= 360) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[6] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,10]
        if ((vga_hcnt >= 361 && vga_hcnt <= 380) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[5] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,11]
        if ((vga_hcnt >= 381 && vga_hcnt <= 400) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[4] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,12]
        if ((vga_hcnt >= 401 && vga_hcnt <= 420) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[3] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,13]
        if ((vga_hcnt >= 421 && vga_hcnt <= 440) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[2] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,14]
        if ((vga_hcnt >= 441 && vga_hcnt <= 460) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[1] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
        
        //[15,15]
        if ((vga_hcnt >= 461 && vga_hcnt <= 480) &&
        	(vga_vcnt >= 381 && vga_vcnt <= 400)) begin
			if(row15[0] == 1'b1)
                begin
                    VGA_R = SCORE_R_ON;
                    VGA_G = SCORE_G_ON;
                    VGA_B = SCORE_B_ON;
                end
            else
                begin
                    VGA_R = SCORE_R_OFF;
                    VGA_G = SCORE_G_OFF;
                    VGA_B = SCORE_B_OFF;
                end
        end
   /************************START BOTTOM ROW***************************************/     
        
                    if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 401) && (vga_vcnt <= 405) ) ) begin
            if(bot_row0[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 406) && (vga_vcnt <= 410) ) ) begin
            if(bot_row1[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 411) && (vga_vcnt <= 415) ) ) begin
            if(bot_row2[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 416) && (vga_vcnt <= 420) ) ) begin
            if(bot_row3[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 421) && (vga_vcnt <= 425) ) ) begin
            if(bot_row4[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 426) && (vga_vcnt <= 430) ) ) begin
            if(bot_row5[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 431) && (vga_vcnt <= 435) ) ) begin
            if(bot_row6[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 436) && (vga_vcnt <= 440) ) ) begin
            if(bot_row7[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 441) && (vga_vcnt <= 445) ) ) begin
            if(bot_row8[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 446) && (vga_vcnt <= 450) ) ) begin
            if(bot_row9[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 451) && (vga_vcnt <= 455) ) ) begin
            if(bot_row10[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 456) && (vga_vcnt <= 460) ) ) begin
            if(bot_row11[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 461) && (vga_vcnt <= 465) ) ) begin
            if(bot_row12[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 466) && (vga_vcnt <= 470) ) ) begin
            if(bot_row13[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 471) && (vga_vcnt <= 475) ) ) begin
            if(bot_row14[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 1) && (vga_hcnt <= 5)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[127] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 6) && (vga_hcnt <= 10)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[126] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 11) && (vga_hcnt <= 15)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[125] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 16) && (vga_hcnt <= 20)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[124] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 21) && (vga_hcnt <= 25)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[123] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 26) && (vga_hcnt <= 30)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[122] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 31) && (vga_hcnt <= 35)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[121] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 36) && (vga_hcnt <= 40)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[120] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 41) && (vga_hcnt <= 45)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[119] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 46) && (vga_hcnt <= 50)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[118] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 51) && (vga_hcnt <= 55)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[117] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 56) && (vga_hcnt <= 60)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[116] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 61) && (vga_hcnt <= 65)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[115] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 66) && (vga_hcnt <= 70)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[114] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 71) && (vga_hcnt <= 75)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[113] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 76) && (vga_hcnt <= 80)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[112] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 81) && (vga_hcnt <= 85)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[111] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 86) && (vga_hcnt <= 90)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[110] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 91) && (vga_hcnt <= 95)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[109] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 96) && (vga_hcnt <= 100)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[108] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 101) && (vga_hcnt <= 105)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[107] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 106) && (vga_hcnt <= 110)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[106] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 111) && (vga_hcnt <= 115)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[105] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 116) && (vga_hcnt <= 120)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[104] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 121) && (vga_hcnt <= 125)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[103] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 126) && (vga_hcnt <= 130)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[102] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 131) && (vga_hcnt <= 135)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[101] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 136) && (vga_hcnt <= 140)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[100] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 141) && (vga_hcnt <= 145)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[99] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 146) && (vga_hcnt <= 150)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[98] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 151) && (vga_hcnt <= 155)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[97] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 156) && (vga_hcnt <= 160)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[96] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 161) && (vga_hcnt <= 165)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[95] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 166) && (vga_hcnt <= 170)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[94] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 171) && (vga_hcnt <= 175)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[93] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 176) && (vga_hcnt <= 180)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[92] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 181) && (vga_hcnt <= 185)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[91] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 186) && (vga_hcnt <= 190)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[90] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 191) && (vga_hcnt <= 195)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[89] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 196) && (vga_hcnt <= 200)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[88] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 201) && (vga_hcnt <= 205)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[87] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 206) && (vga_hcnt <= 210)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[86] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 211) && (vga_hcnt <= 215)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[85] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 216) && (vga_hcnt <= 220)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[84] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 221) && (vga_hcnt <= 225)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[83] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 226) && (vga_hcnt <= 230)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[82] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 231) && (vga_hcnt <= 235)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[81] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 236) && (vga_hcnt <= 240)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[80] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 241) && (vga_hcnt <= 245)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[79] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 246) && (vga_hcnt <= 250)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[78] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 251) && (vga_hcnt <= 255)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[77] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 256) && (vga_hcnt <= 260)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[76] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 261) && (vga_hcnt <= 265)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[75] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 266) && (vga_hcnt <= 270)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[74] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 271) && (vga_hcnt <= 275)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[73] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 276) && (vga_hcnt <= 280)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[72] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 281) && (vga_hcnt <= 285)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[71] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 286) && (vga_hcnt <= 290)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[70] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 291) && (vga_hcnt <= 295)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[69] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 296) && (vga_hcnt <= 300)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[68] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 301) && (vga_hcnt <= 305)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[67] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 306) && (vga_hcnt <= 310)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[66] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 311) && (vga_hcnt <= 315)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[65] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 316) && (vga_hcnt <= 320)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[64] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 321) && (vga_hcnt <= 325)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[63] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 326) && (vga_hcnt <= 330)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[62] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 331) && (vga_hcnt <= 335)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[61] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 336) && (vga_hcnt <= 340)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[60] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 341) && (vga_hcnt <= 345)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[59] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 346) && (vga_hcnt <= 350)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[58] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 351) && (vga_hcnt <= 355)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[57] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 356) && (vga_hcnt <= 360)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[56] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 361) && (vga_hcnt <= 365)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[55] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 366) && (vga_hcnt <= 370)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[54] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 371) && (vga_hcnt <= 375)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[53] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 376) && (vga_hcnt <= 380)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[52] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 381) && (vga_hcnt <= 385)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[51] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 386) && (vga_hcnt <= 390)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[50] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 391) && (vga_hcnt <= 395)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[49] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 396) && (vga_hcnt <= 400)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[48] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 401) && (vga_hcnt <= 405)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[47] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 406) && (vga_hcnt <= 410)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[46] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 411) && (vga_hcnt <= 415)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[45] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 416) && (vga_hcnt <= 420)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[44] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 421) && (vga_hcnt <= 425)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[43] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 426) && (vga_hcnt <= 430)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[42] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 431) && (vga_hcnt <= 435)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[41] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 436) && (vga_hcnt <= 440)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[40] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 441) && (vga_hcnt <= 445)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[39] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 446) && (vga_hcnt <= 450)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[38] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 451) && (vga_hcnt <= 455)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[37] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 456) && (vga_hcnt <= 460)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[36] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 461) && (vga_hcnt <= 465)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[35] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 466) && (vga_hcnt <= 470)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[34] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 471) && (vga_hcnt <= 475)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[33] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 476) && (vga_hcnt <= 480)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[32] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 481) && (vga_hcnt <= 485)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[31] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 486) && (vga_hcnt <= 490)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[30] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 491) && (vga_hcnt <= 495)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[29] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 496) && (vga_hcnt <= 500)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[28] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 501) && (vga_hcnt <= 505)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[27] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 506) && (vga_hcnt <= 510)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[26] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 511) && (vga_hcnt <= 515)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[25] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 516) && (vga_hcnt <= 520)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[24] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 521) && (vga_hcnt <= 525)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[23] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 526) && (vga_hcnt <= 530)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[22] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 531) && (vga_hcnt <= 535)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[21] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 536) && (vga_hcnt <= 540)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[20] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 541) && (vga_hcnt <= 545)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[19] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 546) && (vga_hcnt <= 550)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[18] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 551) && (vga_hcnt <= 555)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[17] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 556) && (vga_hcnt <= 560)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[16] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 561) && (vga_hcnt <= 565)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[15] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 566) && (vga_hcnt <= 570)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[14] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 571) && (vga_hcnt <= 575)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[13] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 576) && (vga_hcnt <= 580)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[12] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 581) && (vga_hcnt <= 585)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[11] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 586) && (vga_hcnt <= 590)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[10] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 591) && (vga_hcnt <= 595)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[9] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 596) && (vga_hcnt <= 600)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[8] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 601) && (vga_hcnt <= 605)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[7] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 606) && (vga_hcnt <= 610)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[6] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 611) && (vga_hcnt <= 615)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[5] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 616) && (vga_hcnt <= 620)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[4] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 621) && (vga_hcnt <= 625)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[3] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 626) && (vga_hcnt <= 630)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[2] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 631) && (vga_hcnt <= 635)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[1] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            
            if ( ( (vga_hcnt >= 636) && (vga_hcnt <= 640)) &&
                ( (vga_vcnt >= 476) && (vga_vcnt <= 480) ) ) begin
            if(bot_row15[0] == 1'b1)
                begin
                    VGA_R = BOT_R_ON;
                    VGA_G = BOT_G_ON;
                    VGA_B = BOT_B_ON;
                end
            else
                begin
                    VGA_R = BOT_R_OFF;
                    VGA_G = BOT_G_OFF;
                    VGA_B = BOT_B_OFF;
                end
            
            end
            

        
    end//else !blank
end

endmodule
